`timescale 1ns / 10ps

module decode(
    input clk,
    input cnd,
    input [3:0] DrA,
    input [3:0] DrB,
    input [63:0] DvalC,
    input [63:0] DvalP,
    input [3:0] Dicode,
    input [3:0] Difun,

    input [3:0] edstE,
    input [3:0] edstM,
    input [3:0] MdstE,
    input [3:0] MdstM,
    input [3:0] WdstE,
    input [3:0] WdstM,

    input [63:0] evalE,
    input [63:0] MvalE,
    input [63:0] mvalM,
    input [63:0] WvalM,
    input [63:0] WvalE,
    
    output reg [63:0] rvalA,
    output reg [63:0] rvalB,

    output reg [63:0] rm0,
    output reg [63:0] rm1,
    output reg [63:0] rm2,
    output reg [63:0] rm3,
    output reg [63:0] rm4,
    output reg [63:0] rm5,
    output reg [63:0] rm6,
    output reg [63:0] rm7,
    output reg [63:0] rm8,
    output reg [63:0] rm9,
    output reg [63:0] rm10,
    output reg [63:0] rm11,
    output reg [63:0] rm12,
    output reg [63:0] rm13,
    output reg [63:0] rm14,

    output reg [63:0] dvalA,
    output reg [63:0] dvalB,
    output reg [63:0] dvalC,
    output reg [3:0] ddstE,
    output reg [3:0] ddstM,
    output reg [3:0] dsrcA,
    output reg [3:0] dsrcB,
    output reg [3:0] dicode,
    output reg [3:0] difun,
    input [3:0] Wicode,
    input [3:0] Wifun,
    input Wcnd
);

reg [63:0]rm[0:14];

initial begin

// ASSIGNED COUNTER VALUES FOR CHECKING OUTPUTS

    rm[0] = 64'd0;
    rm[1] = 64'd1;
    rm[2] = 64'd2;
    rm[3] = 64'd3;
    rm[4] = 64'd4;
    rm[5] = 64'd5;
    rm[6] = 64'd6;
    rm[7] = 64'd7;
    rm[8] = 64'd8;
    rm[9] = 64'd9;
    rm[10] = 64'd10;
    rm[11] = 64'd11;
    rm[12] = 64'd12;
    rm[13] = 64'd13;
    rm[14] = 64'd14;

    rvalA = 64'd0;
    rvalB = 64'd0;
end

// DEFINING PARAMETERS FOR ICODE

parameter HALT = 4'b0000;
parameter NOP = 4'b0001;
parameter CMOVXX = 4'b0010;
parameter IRMOVQ = 4'b0011;
parameter RMMOVQ = 4'b0100;
parameter MRMOVQ = 4'b0101;
parameter OPQ = 4'b0110;
parameter JXX = 4'b0111;
parameter CALL = 4'b1000;
parameter RET = 4'b1001;
parameter PUSHQ = 4'b1010;
parameter POPQ = 4'b1011;

// assigning the intermediates

always @(*)
begin

    case(dicode)

        CMOVXX:
        begin
        dsrcA = DrA;
        ddstE = DrB;
        rvalA = rm[dsrcA];
        end

        IRMOVQ:
        begin
        ddstE = DrB;
        end

        RMMOVQ:
        begin
        dsrcA = DrA;
        dsrcB = DrB;
        rvalA = rm[dsrcA];
        rvalB = rm[dsrcB];
        end

        MRMOVQ:
        begin
        dsrcB = DrB;
        ddstM = DrA;
        rvalB = rm[dsrcB];
        end

        OPQ:
        begin
        dsrcB = DrB;
        dsrcA = DrA;
        ddstE = DrB;
        rvalA = rm[dsrcA];
        rvalB = rm[dsrcB];
        end

        CALL:
        begin
        dsrcB = 4'b0100;
        ddstE = 4'b0100;
        rvalB = rm[4];
        end

        RET:
        begin
        dsrcA = 4'b0100;
        dsrcB = 4'b0100;
        ddstE = 4'b0100;
        rvalA = rm[4];
        rvalB = rm[4];
        end

        PUSHQ:
        begin
        dsrcA = DrA;
        dsrcB = 4'b0100;
        ddstE = 4'b0100;
        rvalA = rm[dsrcA];
        rvalB = rm[4];
        end

        POPQ:
        begin
        dsrcA = 4'b0100;
        dsrcB = 4'b0100;
        ddstE = 4'b0100;
        ddstM = DrA;
        rvalA = rm[4];
        rvalB = rm[4];
        end

    endcase
end

// DATA FORWARDING CASES (REFERED DIRECTLY FROM CLASS SLIDES)

always@(*)
begin
    if(Dicode == JXX || Dicode == CALL)
        dvalA = DvalP;
    else if(dsrcA == edstM)
        dvalA = evalE;
    else if(dsrcA == MdstM)
        dvalA = mvalM;
    else if(dsrcA == MdstE)
        dvalA = MvalE;
    else if(dsrcA == WdstM)
        dvalA = WvalM;
    else if(dsrcA == WdstE)
        dvalA = WvalE;
    else
        dvalA = rvalA;


    if(dsrcB == edstE)
        dvalB = evalE;
    else if(dsrcB == MdstM)
        dvalB = mvalM;
    else if(dsrcB == MdstE)
        dvalB = MvalE;
    else if(dsrcB == WdstM)
        dvalB = WvalM;
    else if(dsrcB == WdstE)
        dvalB = WvalE;
    else
        dvalB = rvalB;
end

// PASSING VALUES FROM INPUT STAGE TO CURRENT STAGE

always@(*)
begin
    dicode = Dicode;
    difun = Difun;
    dvalC = DvalC;
end

// WRITE BACK IS WRITTEN INSIDE DECODE CUZ OUR CODE WAS NOT ALLOWING TO CHANGE VALUES OF REGISTERS WHICH WERE DECLARED AS WIRES IN THE PROCPIPE SO WE HAD TO DEFINE A SINGLE MODULE WITH THOSE REGISTERS AS OUTPUTS SO THAT WE CAN CHANGE THEM ONCE AND FOR ALL HERE ONLY

always @ (negedge clk)
    begin
        if(Wicode == CMOVXX && Wifun == 4'b0)
        begin
            rm[WdstE] = WvalE;
        end
        if(Wicode == CMOVXX && Wifun != 4'b0 && Wcnd == 1)
        begin
            // if(cnd)
            // begin
                 rm[WdstE] = WvalE;
            // end
            // else
            // begin
            //     rm[14] = valE;
            // end

            // UGHHHHHHH SILLY ERRORRRRRRRRRRRRR!!!!!!!!!!!!!!

            // case(cnd)

            // 1'b1:
            // begin
            //     rm[rB] = valE;
            // end

            // default:
            // begin
            //     rm[14] = valE;
            // end

            // endcase
        end

        else if(Wicode == IRMOVQ)
        begin
        rm[WdstE] = WvalE;
        // rm[4] = 5; // FOR TESTING PURPOSES ONLY
        end

        else if(Wicode == MRMOVQ)
        begin
        rm[WdstM] = WvalM;
        end

        else if(Wicode == OPQ)
        begin
        rm[WdstE] = WvalE;
        end

        else if(Wicode == CALL)
        begin
        rm[4] = WvalE;
        end

        else if(Wicode == RET)
        begin
        rm[4] = WvalE;
        end

        else if(Wicode == PUSHQ)
        begin
        rm[4] = WvalE;
        end

        else if(Wicode == POPQ)
        begin
        rm[4] = WvalE;
        rm[WdstM] = WvalM;
        end

        // ASSIGNING REG VARIABLES TO SEE OUTPUTS AS ARRAY ELEMENTS $MONITOR WAS NOT SUPPORTING

        rm0 = rm[0];
        rm1 = rm[1];
        rm2 = rm[2];
        rm3 = rm[3];
        rm4 = rm[4];
        rm5 = rm[5];
        rm6 = rm[6];
        rm7 = rm[7];
        rm8 = rm[8];
        rm9 = rm[9];
        rm10 = rm[10];
        rm11 = rm[11];
        rm12 = rm[12];
        rm13 = rm[13];
        rm14 = rm[14];

end

endmodule



   

