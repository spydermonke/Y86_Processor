`timescale 1ns / 1ps

module andg(p,q,r);

input p;
input q;
output r;

and gate1(r,p,q);

endmodule